library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity IMemory_16_16 is
	generic(N        : integer := 16);
	port(Enable      : in  std_logic;
		  registAdress: in  std_logic_vector(N-1 downto 0);
		  readData    : out std_logic_vector(N-1 downto 0));
end IMemory_16_16;

architecture Behavioral of IMemory_16_16 is
	subtype TDataWord is std_logic_vector(N-1 downto 0);
	type TROM is array (0 to N-1) of TDataWord;
	constant c_memory: TROM := ("0110000010000000", "1000000100000001", "0010010100110110", "0010000111000000",
										 "1000100100000001", "0010010100110110", "0011000111000000", "1000100100000001", 
										 "0010010100110110", "0011000111000000", "1100000100000010", "1100001000000011");
	begin
		if(Enable <= '1') then
			readData <= c_memory(to_integer(unsigned(registAdress)));
		end if;
end Behavioral;